module pc1(input [1:64]key, output [1:56]key_pc1);
assign key_pc1[1] = key[57];
assign key_pc1[2] = key[49];
assign key_pc1[3] = key[41];
assign key_pc1[4] = key[33];
assign key_pc1[5] = key[25];
assign key_pc1[6] = key[17];
assign key_pc1[7] = key[9];
assign key_pc1[8] = key[1];
assign key_pc1[9] = key[58];
assign key_pc1[10] = key[50];
assign key_pc1[11] = key[42];
assign key_pc1[12] = key[34];
assign key_pc1[13] = key[26];
assign key_pc1[14] = key[18];
assign key_pc1[15] = key[10];
assign key_pc1[16] = key[2];
assign key_pc1[17] = key[59];
assign key_pc1[18] = key[51];
assign key_pc1[19] = key[43];
assign key_pc1[20] = key[35];
assign key_pc1[21] = key[27];
assign key_pc1[22] = key[19];
assign key_pc1[23] = key[11];
assign key_pc1[24] = key[3];
assign key_pc1[25] = key[60];
assign key_pc1[26] = key[52];
assign key_pc1[27] = key[44];
assign key_pc1[28] = key[36];
assign key_pc1[29] = key[63];
assign key_pc1[30] = key[55];
assign key_pc1[31] = key[47];
assign key_pc1[32] = key[39];
assign key_pc1[33] = key[31];
assign key_pc1[34] = key[23];
assign key_pc1[35] = key[15];
assign key_pc1[36] = key[7];
assign key_pc1[37] = key[62];
assign key_pc1[38] = key[54];
assign key_pc1[39] = key[46];
assign key_pc1[40] = key[38];
assign key_pc1[41] = key[30];
assign key_pc1[42] = key[22];
assign key_pc1[43] = key[14];
assign key_pc1[44] = key[6];
assign key_pc1[45] = key[61];
assign key_pc1[46] = key[53];
assign key_pc1[47] = key[45];
assign key_pc1[48] = key[37];
assign key_pc1[49] = key[29];
assign key_pc1[50] = key[21];
assign key_pc1[51] = key[13];
assign key_pc1[52] = key[5];
assign key_pc1[53] = key[28];
assign key_pc1[54] = key[20];
assign key_pc1[55] = key[12];
assign key_pc1[56] = key[4];
endmodule